// ============================================================================
// Module: cpu_top
// Author: Zhong Litao
// Created: 2025-09-25
// Description: 
// top connection
// ============================================================================

`timescale 1ns / 1ps
import my_pkg.sv::*;
module cpu_top
(
    input wire         clk      ,
    input wire         rst_n    
);


endmodule